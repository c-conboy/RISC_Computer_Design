module ror(output[31:0]C, input[31:0]A);
	assign C[31] = A[0];
	assign C[30:0] = A[31:1];
endmodule
	